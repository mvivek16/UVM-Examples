`timescale 1ns/10ps

package mypackage;
	integer a;
endpackage
