`include "_40_cat_dog_pkg.sv"

import uvm_pkg::*;
import cat_dog::*;
//`include "uvm_macros.svh"

module top;
	initial
		run_test();
endmodule
